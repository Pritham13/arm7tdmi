module Control (
    input
);
    
endmodule