module ALU_decoder (
    input opcode
);
    
endmodule